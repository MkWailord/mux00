entity fa00 is
port(
	C00: in std_logic;
	A00: in std_logic;
	B00: in std_logic;
	S00: out std_logic;
	C01: out std_logic
);
end fa00;

architecture fa0 